
  module InlineBlackBoxLut(
      input  [7:0] rom_addr,
      output [7:0] rom_dout
      );
   wire [7:0] rom_256_8 [0:255];  // 256 words in total
   assign rom_dout = {1'b1,rom_256_8[rom_addr]};
   assign rom_256_8[0] = 7 'b1111111;
   assign rom_256_8[1] = 7 'b1111110;
   assign rom_256_8[2] = 7 'b1111101;
   assign rom_256_8[3] = 7 'b1111100;
   assign rom_256_8[4] = 7 'b1111011;
   assign rom_256_8[5] = 7 'b1111010;
   assign rom_256_8[6] = 7 'b1111001;
   assign rom_256_8[7] = 7 'b1111000;
   assign rom_256_8[8] = 7 'b1110111;
   assign rom_256_8[9] = 7 'b1110110;
   assign rom_256_8[10] = 7 'b1110101;
   assign rom_256_8[11] = 7 'b1110100;
   assign rom_256_8[12] = 7 'b1110011;
   assign rom_256_8[13] = 7 'b1110011;
   assign rom_256_8[14] = 7 'b1110010;
   assign rom_256_8[15] = 7 'b1110001;
   assign rom_256_8[16] = 7 'b1110000;
   assign rom_256_8[17] = 7 'b1101111;
   assign rom_256_8[18] = 7 'b1101110;
   assign rom_256_8[19] = 7 'b1101101;
   assign rom_256_8[20] = 7 'b1101100;
   assign rom_256_8[21] = 7 'b1101100;
   assign rom_256_8[22] = 7 'b1101011;
   assign rom_256_8[23] = 7 'b1101010;
   assign rom_256_8[24] = 7 'b1101001;
   assign rom_256_8[25] = 7 'b1101000;
   assign rom_256_8[26] = 7 'b1101000;
   assign rom_256_8[27] = 7 'b1100111;
   assign rom_256_8[28] = 7 'b1100110;
   assign rom_256_8[29] = 7 'b1100101;
   assign rom_256_8[30] = 7 'b1100100;
   assign rom_256_8[31] = 7 'b1100100;
   assign rom_256_8[32] = 7 'b1100011;
   assign rom_256_8[33] = 7 'b1100010;
   assign rom_256_8[34] = 7 'b1100001;
   assign rom_256_8[35] = 7 'b1100000;
   assign rom_256_8[36] = 7 'b1100000;
   assign rom_256_8[37] = 7 'b1011111;
   assign rom_256_8[38] = 7 'b1011110;
   assign rom_256_8[39] = 7 'b1011101;
   assign rom_256_8[40] = 7 'b1011101;
   assign rom_256_8[41] = 7 'b1011100;
   assign rom_256_8[42] = 7 'b1011011;
   assign rom_256_8[43] = 7 'b1011010;
   assign rom_256_8[44] = 7 'b1011010;
   assign rom_256_8[45] = 7 'b1011001;
   assign rom_256_8[46] = 7 'b1011000;
   assign rom_256_8[47] = 7 'b1011000;
   assign rom_256_8[48] = 7 'b1010111;
   assign rom_256_8[49] = 7 'b1010110;
   assign rom_256_8[50] = 7 'b1010110;
   assign rom_256_8[51] = 7 'b1010101;
   assign rom_256_8[52] = 7 'b1010100;
   assign rom_256_8[53] = 7 'b1010011;
   assign rom_256_8[54] = 7 'b1010011;
   assign rom_256_8[55] = 7 'b1010010;
   assign rom_256_8[56] = 7 'b1010001;
   assign rom_256_8[57] = 7 'b1010001;
   assign rom_256_8[58] = 7 'b1010000;
   assign rom_256_8[59] = 7 'b1001111;
   assign rom_256_8[60] = 7 'b1001111;
   assign rom_256_8[61] = 7 'b1001110;
   assign rom_256_8[62] = 7 'b1001110;
   assign rom_256_8[63] = 7 'b1001101;
   assign rom_256_8[64] = 7 'b1001100;
   assign rom_256_8[65] = 7 'b1001100;
   assign rom_256_8[66] = 7 'b1001011;
   assign rom_256_8[67] = 7 'b1001010;
   assign rom_256_8[68] = 7 'b1001010;
   assign rom_256_8[69] = 7 'b1001001;
   assign rom_256_8[70] = 7 'b1001000;
   assign rom_256_8[71] = 7 'b1001000;
   assign rom_256_8[72] = 7 'b1000111;
   assign rom_256_8[73] = 7 'b1000111;
   assign rom_256_8[74] = 7 'b1000110;
   assign rom_256_8[75] = 7 'b1000101;
   assign rom_256_8[76] = 7 'b1000101;
   assign rom_256_8[77] = 7 'b1000100;
   assign rom_256_8[78] = 7 'b1000100;
   assign rom_256_8[79] = 7 'b1000011;
   assign rom_256_8[80] = 7 'b1000011;
   assign rom_256_8[81] = 7 'b1000010;
   assign rom_256_8[82] = 7 'b1000001;
   assign rom_256_8[83] = 7 'b1000001;
   assign rom_256_8[84] = 7 'b1000000;
   assign rom_256_8[85] = 7 'b1000000;
   assign rom_256_8[86] = 7 'b0111111;
   assign rom_256_8[87] = 7 'b0111111;
   assign rom_256_8[88] = 7 'b0111110;
   assign rom_256_8[89] = 7 'b0111101;
   assign rom_256_8[90] = 7 'b0111101;
   assign rom_256_8[91] = 7 'b0111100;
   assign rom_256_8[92] = 7 'b0111100;
   assign rom_256_8[93] = 7 'b0111011;
   assign rom_256_8[94] = 7 'b0111011;
   assign rom_256_8[95] = 7 'b0111010;
   assign rom_256_8[96] = 7 'b0111010;
   assign rom_256_8[97] = 7 'b0111001;
   assign rom_256_8[98] = 7 'b0111001;
   assign rom_256_8[99] = 7 'b0111000;
   assign rom_256_8[100] = 7 'b0111000;
   assign rom_256_8[101] = 7 'b0110111;
   assign rom_256_8[102] = 7 'b0110111;
   assign rom_256_8[103] = 7 'b0110110;
   assign rom_256_8[104] = 7 'b0110110;
   assign rom_256_8[105] = 7 'b0110101;
   assign rom_256_8[106] = 7 'b0110101;
   assign rom_256_8[107] = 7 'b0110100;
   assign rom_256_8[108] = 7 'b0110100;
   assign rom_256_8[109] = 7 'b0110011;
   assign rom_256_8[110] = 7 'b0110011;
   assign rom_256_8[111] = 7 'b0110010;
   assign rom_256_8[112] = 7 'b0110010;
   assign rom_256_8[113] = 7 'b0110001;
   assign rom_256_8[114] = 7 'b0110001;
   assign rom_256_8[115] = 7 'b0110000;
   assign rom_256_8[116] = 7 'b0110000;
   assign rom_256_8[117] = 7 'b0101111;
   assign rom_256_8[118] = 7 'b0101111;
   assign rom_256_8[119] = 7 'b0101110;
   assign rom_256_8[120] = 7 'b0101110;
   assign rom_256_8[121] = 7 'b0101101;
   assign rom_256_8[122] = 7 'b0101101;
   assign rom_256_8[123] = 7 'b0101100;
   assign rom_256_8[124] = 7 'b0101100;
   assign rom_256_8[125] = 7 'b0101100;
   assign rom_256_8[126] = 7 'b0101011;
   assign rom_256_8[127] = 7 'b0101011;
   assign rom_256_8[128] = 7 'b0101010;
   assign rom_256_8[129] = 7 'b0101010;
   assign rom_256_8[130] = 7 'b0101001;
   assign rom_256_8[131] = 7 'b0101001;
   assign rom_256_8[132] = 7 'b0101000;
   assign rom_256_8[133] = 7 'b0101000;
   assign rom_256_8[134] = 7 'b0101000;
   assign rom_256_8[135] = 7 'b0100111;
   assign rom_256_8[136] = 7 'b0100111;
   assign rom_256_8[137] = 7 'b0100110;
   assign rom_256_8[138] = 7 'b0100110;
   assign rom_256_8[139] = 7 'b0100101;
   assign rom_256_8[140] = 7 'b0100101;
   assign rom_256_8[141] = 7 'b0100101;
   assign rom_256_8[142] = 7 'b0100100;
   assign rom_256_8[143] = 7 'b0100100;
   assign rom_256_8[144] = 7 'b0100011;
   assign rom_256_8[145] = 7 'b0100011;
   assign rom_256_8[146] = 7 'b0100011;
   assign rom_256_8[147] = 7 'b0100010;
   assign rom_256_8[148] = 7 'b0100010;
   assign rom_256_8[149] = 7 'b0100001;
   assign rom_256_8[150] = 7 'b0100001;
   assign rom_256_8[151] = 7 'b0100001;
   assign rom_256_8[152] = 7 'b0100000;
   assign rom_256_8[153] = 7 'b0100000;
   assign rom_256_8[154] = 7 'b0011111;
   assign rom_256_8[155] = 7 'b0011111;
   assign rom_256_8[156] = 7 'b0011111;
   assign rom_256_8[157] = 7 'b0011110;
   assign rom_256_8[158] = 7 'b0011110;
   assign rom_256_8[159] = 7 'b0011101;
   assign rom_256_8[160] = 7 'b0011101;
   assign rom_256_8[161] = 7 'b0011101;
   assign rom_256_8[162] = 7 'b0011100;
   assign rom_256_8[163] = 7 'b0011100;
   assign rom_256_8[164] = 7 'b0011100;
   assign rom_256_8[165] = 7 'b0011011;
   assign rom_256_8[166] = 7 'b0011011;
   assign rom_256_8[167] = 7 'b0011010;
   assign rom_256_8[168] = 7 'b0011010;
   assign rom_256_8[169] = 7 'b0011010;
   assign rom_256_8[170] = 7 'b0011001;
   assign rom_256_8[171] = 7 'b0011001;
   assign rom_256_8[172] = 7 'b0011001;
   assign rom_256_8[173] = 7 'b0011000;
   assign rom_256_8[174] = 7 'b0011000;
   assign rom_256_8[175] = 7 'b0011000;
   assign rom_256_8[176] = 7 'b0010111;
   assign rom_256_8[177] = 7 'b0010111;
   assign rom_256_8[178] = 7 'b0010111;
   assign rom_256_8[179] = 7 'b0010110;
   assign rom_256_8[180] = 7 'b0010110;
   assign rom_256_8[181] = 7 'b0010101;
   assign rom_256_8[182] = 7 'b0010101;
   assign rom_256_8[183] = 7 'b0010101;
   assign rom_256_8[184] = 7 'b0010100;
   assign rom_256_8[185] = 7 'b0010100;
   assign rom_256_8[186] = 7 'b0010100;
   assign rom_256_8[187] = 7 'b0010011;
   assign rom_256_8[188] = 7 'b0010011;
   assign rom_256_8[189] = 7 'b0010011;
   assign rom_256_8[190] = 7 'b0010010;
   assign rom_256_8[191] = 7 'b0010010;
   assign rom_256_8[192] = 7 'b0010010;
   assign rom_256_8[193] = 7 'b0010001;
   assign rom_256_8[194] = 7 'b0010001;
   assign rom_256_8[195] = 7 'b0010001;
   assign rom_256_8[196] = 7 'b0010000;
   assign rom_256_8[197] = 7 'b0010000;
   assign rom_256_8[198] = 7 'b0010000;
   assign rom_256_8[199] = 7 'b0010000;
   assign rom_256_8[200] = 7 'b0001111;
   assign rom_256_8[201] = 7 'b0001111;
   assign rom_256_8[202] = 7 'b0001111;
   assign rom_256_8[203] = 7 'b0001110;
   assign rom_256_8[204] = 7 'b0001110;
   assign rom_256_8[205] = 7 'b0001110;
   assign rom_256_8[206] = 7 'b0001101;
   assign rom_256_8[207] = 7 'b0001101;
   assign rom_256_8[208] = 7 'b0001101;
   assign rom_256_8[209] = 7 'b0001100;
   assign rom_256_8[210] = 7 'b0001100;
   assign rom_256_8[211] = 7 'b0001100;
   assign rom_256_8[212] = 7 'b0001100;
   assign rom_256_8[213] = 7 'b0001011;
   assign rom_256_8[214] = 7 'b0001011;
   assign rom_256_8[215] = 7 'b0001011;
   assign rom_256_8[216] = 7 'b0001010;
   assign rom_256_8[217] = 7 'b0001010;
   assign rom_256_8[218] = 7 'b0001010;
   assign rom_256_8[219] = 7 'b0001001;
   assign rom_256_8[220] = 7 'b0001001;
   assign rom_256_8[221] = 7 'b0001001;
   assign rom_256_8[222] = 7 'b0001001;
   assign rom_256_8[223] = 7 'b0001000;
   assign rom_256_8[224] = 7 'b0001000;
   assign rom_256_8[225] = 7 'b0001000;
   assign rom_256_8[226] = 7 'b0000111;
   assign rom_256_8[227] = 7 'b0000111;
   assign rom_256_8[228] = 7 'b0000111;
   assign rom_256_8[229] = 7 'b0000111;
   assign rom_256_8[230] = 7 'b0000110;
   assign rom_256_8[231] = 7 'b0000110;
   assign rom_256_8[232] = 7 'b0000110;
   assign rom_256_8[233] = 7 'b0000110;
   assign rom_256_8[234] = 7 'b0000101;
   assign rom_256_8[235] = 7 'b0000101;
   assign rom_256_8[236] = 7 'b0000101;
   assign rom_256_8[237] = 7 'b0000100;
   assign rom_256_8[238] = 7 'b0000100;
   assign rom_256_8[239] = 7 'b0000100;
   assign rom_256_8[240] = 7 'b0000100;
   assign rom_256_8[241] = 7 'b0000011;
   assign rom_256_8[242] = 7 'b0000011;
   assign rom_256_8[243] = 7 'b0000011;
   assign rom_256_8[244] = 7 'b0000011;
   assign rom_256_8[245] = 7 'b0000010;
   assign rom_256_8[246] = 7 'b0000010;
   assign rom_256_8[247] = 7 'b0000010;
   assign rom_256_8[248] = 7 'b0000010;
   assign rom_256_8[249] = 7 'b0000001;
   assign rom_256_8[250] = 7 'b0000001;
   assign rom_256_8[251] = 7 'b0000001;
   assign rom_256_8[252] = 7 'b0000001;
   assign rom_256_8[253] = 7 'b0000000;
   assign rom_256_8[254] = 7 'b0000000;
   assign rom_256_8[255] = 7 'b0000000;
   endmodule
   